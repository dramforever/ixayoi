typedef Bit#(32)    Word;
typedef Bit#(4)     BStrb;

typedef Bit#(32)    Instr;
typedef Bit#(5)     RegNum;
typedef Bit#(7)     Opcode;
typedef Bit#(7)     Funct7;
typedef Bit#(3)     Funct3;

typedef Int#(32)    SWord;
